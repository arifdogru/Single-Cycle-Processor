module mips_ALU_32Bit_MSB();

endmodule