module shiftLeft(inp,result);

input [31:0] inp;
output [31:0] result;

assign result = inp <<2; 

endmodule